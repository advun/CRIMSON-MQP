`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/31/2025 02:41:42 PM
// Design Name: 
// Module Name: SARADC
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SARADC(
    input clk,
    input start,
    input reset_n,
    output [9:0] D,
    output [9:0] bitctrl
    );
    
    
endmodule
